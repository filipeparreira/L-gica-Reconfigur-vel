library verilog;
use verilog.vl_types.all;
entity Atividade1_vlg_vec_tst is
end Atividade1_vlg_vec_tst;
