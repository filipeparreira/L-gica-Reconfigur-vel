library ieee;
use ieee.std_logic_1164;

entity atividade7 is port(
	reset, pause, mudar, up, down: in std_logic;
	ssd1, ssd2, ssd3, ssd4: out std_logic_vector(6 DOWNTO 0)
);
end atividade7;

architecture main of atividade7 is 

begin 



end main;