library verilog;
use verilog.vl_types.all;
entity atividade_2_vlg_vec_tst is
end atividade_2_vlg_vec_tst;
