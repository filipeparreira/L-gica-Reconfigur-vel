library verilog;
use verilog.vl_types.all;
entity atividade_2_vlg_check_tst is
    port(
        sirene          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end atividade_2_vlg_check_tst;
