library verilog;
use verilog.vl_types.all;
entity atividade_2_vlg_sample_tst is
    port(
        c               : in     vl_logic;
        f               : in     vl_logic;
        m               : in     vl_logic;
        p               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end atividade_2_vlg_sample_tst;
