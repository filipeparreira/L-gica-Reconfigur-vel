library verilog;
use verilog.vl_types.all;
entity atividade_2 is
    port(
        p               : in     vl_logic;
        m               : in     vl_logic;
        f               : in     vl_logic;
        c               : in     vl_logic;
        sirene          : out    vl_logic
    );
end atividade_2;
