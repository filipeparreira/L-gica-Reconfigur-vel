library verilog;
use verilog.vl_types.all;
entity atividade_4_vlg_vec_tst is
end atividade_4_vlg_vec_tst;
