library verilog;
use verilog.vl_types.all;
entity atividade_4_vlg_check_tst is
    port(
        saida           : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end atividade_4_vlg_check_tst;
