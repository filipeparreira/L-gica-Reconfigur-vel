library ieee;
use ieee.std_logic_1164;

package ssd is 
	procedure ssd_numbers(in1, in2, in3, in4: in std_logic_vector(6 downto 0);
									out1, out2, out3, out4: out std_logic_vector(6 downto 0));
end ssd;

package body ssd is
	procedure ssd_numbers(in1, in2, in3, in4: in std_logic_vector(6 downto 0);
									out1, out2, out3, out4: out std_logic_vector(6 downto 0)) is 
	begin 
	
	end ssd_numbers;
end ssd;